`timescale 1ns / 1ps
//
// WIDTH: bits in register hdata & vdata
// HSIZE: horizontal size of visible field 
// HFP: horizontal front of pulse
// HSP: horizontal stop of pulse
// HMAX: horizontal max size of value
// VSIZE: vertical size of visible field 
// VFP: vertical front of pulse
// VSP: vertical stop of pulse
// VMAX: vertical max size of value
// HSPP: horizontal synchro pulse polarity (0 - negative, 1 - positive)
// VSPP: vertical synchro pulse polarity (0 - negative, 1 - positive)
//
module video
#(parameter WIDTH = 0, HSIZE = 0, HFP = 0, HSP = 0, HMAX = 0, VSIZE = 0, VFP = 0, VSP = 0, VMAX = 0, HSPP = 0, VSPP = 0)
(
    input wire clk,
    input wire rst_n,
    output wire hsync,
    output wire vsync,
    output reg [WIDTH - 1:0] hdata,
    output reg [WIDTH - 1:0] vdata
);

//    initial begin
//        hdata = 'b0;
//        vdata = 'b0;
//    end
    
//    always_ff@(posedge clk)begin
//        if(rst_n)begin
//            hdata<=0;
//            vdata<=0;
//        end
//    end
    
    always_ff@(posedge clk)begin
        if(rst_n)begin
            hdata<=0;
            vdata<=0;
        end
        else begin
            if (hdata == (HMAX - 1))begin
                hdata <= 0;
                if (vdata == (VMAX - 1))
                    vdata <= 0;
                else
                    vdata <= vdata + 1;
            end
            else begin
                hdata <= hdata + 1;
            end
        end
    end
    
    // hdata
//    always @ (posedge clk)
//    begin
//        if (hdata == (HMAX - 1))
//            hdata <= 0;
//        else
//            hdata <= hdata + 1;
//    end

//    // vdata
//    always @ (posedge clk)
//    begin
//        if (hdata == (HMAX - 1)) 
//        begin
//            if (vdata == (VMAX - 1))
//                vdata <= 0;
//            else
//                vdata <= vdata + 1;
//        end
//    end

    // hsync & vsync & blank
    assign hsync = ((hdata >= HFP) && (hdata < HSP)) ? HSPP : !HSPP;
    assign vsync = ((vdata >= VFP) && (vdata < VSP)) ? VSPP : !VSPP;
//    assign data_enable = ((hdata < HSIZE) & (vdata < VSIZE));

endmodule
